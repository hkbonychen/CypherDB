library verilog;
use verilog.vl_types.all;
entity or1200_ctrl is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        except_flushpipe: in     vl_logic;
        extend_flush    : in     vl_logic;
        if_flushpipe    : out    vl_logic;
        id_flushpipe    : out    vl_logic;
        ex_flushpipe    : out    vl_logic;
        wb_flushpipe    : out    vl_logic;
        id_freeze       : in     vl_logic;
        ex_freeze       : in     vl_logic;
        wb_freeze       : in     vl_logic;
        if_insn         : in     vl_logic_vector(31 downto 0);
        id_insn         : out    vl_logic_vector(31 downto 0);
        ex_insn         : out    vl_logic_vector(31 downto 0);
        abort_mvspr     : in     vl_logic;
        id_branch_op    : out    vl_logic_vector(2 downto 0);
        ex_branch_op    : out    vl_logic_vector(2 downto 0);
        ex_branch_taken : in     vl_logic;
        pc_we           : in     vl_logic;
        rf_addra        : out    vl_logic_vector(4 downto 0);
        rf_addrb        : out    vl_logic_vector(4 downto 0);
        rf_rda          : out    vl_logic;
        rf_rdb          : out    vl_logic;
        alu_op          : out    vl_logic_vector(4 downto 0);
        alu_op2         : out    vl_logic_vector(3 downto 0);
        mac_op          : out    vl_logic_vector(2 downto 0);
        comp_op         : out    vl_logic_vector(3 downto 0);
        rf_addrw        : out    vl_logic_vector(4 downto 0);
        rfwb_op         : out    vl_logic_vector(3 downto 0);
        fpu_op          : out    vl_logic_vector(7 downto 0);
        wb_insn         : out    vl_logic_vector(31 downto 0);
        id_simm         : out    vl_logic_vector(31 downto 0);
        ex_simm         : out    vl_logic_vector(31 downto 0);
        id_branch_addrtarget: out    vl_logic_vector(31 downto 2);
        ex_branch_addrtarget: out    vl_logic_vector(31 downto 2);
        sel_a           : out    vl_logic_vector(1 downto 0);
        sel_b           : out    vl_logic_vector(1 downto 0);
        id_lsu_op       : out    vl_logic_vector(3 downto 0);
        cust5_op        : out    vl_logic_vector(4 downto 0);
        cust5_limm      : out    vl_logic_vector(5 downto 0);
        id_pc           : in     vl_logic_vector(31 downto 0);
        ex_pc           : in     vl_logic_vector(31 downto 0);
        du_hwbkpt       : in     vl_logic;
        multicycle      : out    vl_logic_vector(2 downto 0);
        wait_on         : out    vl_logic_vector(1 downto 0);
        wbforw_valid    : in     vl_logic;
        sig_syscall     : out    vl_logic;
        sig_trap        : out    vl_logic;
        force_dslot_fetch: out    vl_logic;
        no_more_dslot   : out    vl_logic;
        id_void         : out    vl_logic;
        ex_void         : out    vl_logic;
        ex_spr_read     : out    vl_logic;
        ex_spr_write    : out    vl_logic;
        id_mac_op       : out    vl_logic_vector(2 downto 0);
        id_macrc_op     : out    vl_logic;
        ex_macrc_op     : out    vl_logic;
        rfe             : out    vl_logic;
        except_illegal  : out    vl_logic;
        dc_no_writethrough: out    vl_logic
    );
end or1200_ctrl;
