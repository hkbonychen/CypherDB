library verilog;
use verilog.vl_types.all;
entity or1200_iwb_biu is
end or1200_iwb_biu;
